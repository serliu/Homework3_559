module FSM_CRC_checker();



endmodule 